
module EX_MEM(reset,clk,JumpPC_in,JumpPC_out,zero_in,zero_out);

input reset, clk; 
input[31:0] JumpPC_in;
output[31:0] JumpPC_out; 



endmodule 