
module shift3 (in, out);

input [127:0] in;
output [127:0] out;

assign out = in<<3; 


endmodule 
