
module IF_ID (PC_adderOut,instruction1,instruction2,