
module Execute (readDataRA_EX, readDataRB_EX, readDataRC_EX, opcode_EX,
	        imm7, imm10, imm16, imm18, 
		result_EX, latency_EX, branch_PC, branch_flag,local_store_address);

                          

//Jump Branch datapath 
input signed [127:0] readDataRA_EX; 
input signed [127:0] readDataRB_EX;
input signed [127:0] readDataRC_EX;
input [6:0] opcode_EX;  
input signed [6:0] imm7; 
input signed [9:0] imm10;
input signed [15:0] imm16;
input signed  [17:0] imm18;

output logic [31:0] branch_PC,local_store_address; //new PC address
logic [17:0] branch_PC_p1; //add first two bits to PC address 
logic [31:0] branch_PC_p2; 
logic [7:0] temp_b,temp_c; // 8 bit temp number 		   
logic [31:0] temp_bbbb;
logic [15:0] temp_r,temp_s,temp_k;	

output [127:0] result_EX; //perhaps not needed, if we have 
output logic [2:0] latency_EX; 
output logic branch_flag=0;	//set default to 0
logic [127:0] RT;
logic [127:0] RA;
logic [127:0] RB; 
logic [127:0] RC;
logic [127:0] unsigned_RA;
logic [127:0] unsigned_RB;
logic [127:0] unsigned_RC;	
shortreal float_RA;
shortreal float_RB;
shortreal float_RC; 

logic [15:0] imm_extended;
logic [31:0] imm_extended_32; 
logic [31:0] temp_32,temp_u,temp_t,temp_t1,temp_t2,temp_t3;  
logic [15:0] unsigned_imm_extended;
logic [31:0] unsigned_imm_extended_32;

assign result_EX     = RT; 
assign RA = readDataRA_EX; 
assign RB = readDataRB_EX; 
assign RC = readDataRC_EX; 

assign unsigned_RA= unsigned'(RA);

assign unsigned_RB= unsigned'(RB);

assign unsigned_RC= unsigned'(RC);	 
assign float_RA= shortreal'(RA); 

assign float_RB= shortreal'(RB);
assign float_RC= shortreal'(RC);

assign branch_PC_p1={imm16,{2{1'b0}}}; 	//add two extra bits 
assign branch_PC_p2={{14{branch_PC_p1[17]}},branch_PC_p1}; 
//assign branch_PC=branch_PC_p2&32'hFFFFFFFC; //extend to 32 bits  
//assign unsigned_imm_extended=unsigned'(imm_extended);  
//assign unsigned_imm_extended_32=unsigned'(imm_extended_32);


always_comb begin
	case(opcode_EX) 
		7'd5: begin //add halfword 
			latency_EX= 3-1; 
			RT[0+:16] = RA[0+:16]+RB[0+:16]; //bytes 0 and 1
			RT[16+:16]=RA[16+:16]+RB[16+:16]; //bytes 2 and 3
			RT[32+:16]=RA[32+:16]+RB[32+:16]; //bytes 4 and 5
			RT[48+:16]=RA[48+:16]+RB[48+:16]; //bytes 6 and 7
			RT[64+:16]=RA[64+:16]+RB[64+:16]; //bytes 8 and 9 
			RT[80+:16]=RA[80+:16]+RB[80+:16]; //bytes 10 and 11 
			RT[96+:16]=RA[96+:16]+RB[96+:16]; //bytes 12 and 13
			RT[112+:16]=RA[112+:16]+RB[112+:16]; //bytes 14 and 15 

		end 
		
	7'd6: //add	halfword immediate 
	begin 
	        latency_EX= 3-1; 	 //add halfword immediate
			imm_extended={ {6{imm10[9]}},imm10};
			RT[0+:16] = RA[0+:16]+imm_extended;
			RT[16+:16]=RA[16+:16]+imm_extended;
			RT[32+:16]=RA[32+:16]+imm_extended;
			RT[48+:16]=RA[48+:16]+imm_extended;
			RT[64+:16]=RA[64+:16]+imm_extended;
			RT[80+:16]=RA[80+:16]+imm_extended;
			RT[96+:16]=RA[96+:16]+imm_extended;
			RT[112+:16]=RA[112+:16]+imm_extended; 
	end 
	7'd7: //add word 
	begin 
	        RT[0+:32] = RA[0+:32]+RB[0+:32]; //bytes 0 and 3
			RT[32+:32]=RA[32+:32]+RB[32+:32]; //bytes 4 and 7
			RT[64+:32]=RA[64+:32]+RB[64+:32]; //bytes 8 and 11
			RT[96+:32]=RA[96+:32]+RB[96+:32]; //bytes 12 and 15
				
		
		
		
	end   
	7'd8:
	begin 
	        latency_EX= 3-1; //add word immediate	   
	 		imm_extended_32={ {22{imm10[9]}},imm10};
			RT[0+:32] = RA[0+:32]+imm_extended_32;
			RT[32+:32]=RA[32+:32]+imm_extended_32;
			RT[64+:32]=RA[64+:32]+imm_extended_32;
			RT[96+:32]=RA[96+:32]+imm_extended_32; 
			
		
		
	end	 
	7'd9: 
	begin  //subtract from halfword 
	        latency_EX= 3-1;  
			RT[0+:16] = RB[0+:16]+ (~RA[0+:16]+1); //bytes 0 and 1
			RT[16+:16]=RB[16+:16]+(~RA[16+:16]+1); //bytes 2 and 3
			RT[32+:16]=RB[32+:16]+(~RA[32+:16]+1); //bytes 4 and 5
			RT[48+:16]=RB[48+:16]+(~RA[48+:16]+1); //bytes 6 and 7
			RT[64+:16]=RB[64+:16]+(~RA[64+:16]+1); //bytes 8 and 9 
			RT[80+:16]=RB[80+:16]+(~RA[80+:16]+1); //bytes 10 and 11 
			RT[96+:16]=RB[96+:16]+(~RA[96+:16]+1); //bytes 12 and 13
			RT[112+:16]=RB[112+:16]+(~RA[112+:16]+1); //bytes 14 and 15 	
		
		
	end
	7'd10: begin	 //subtract from halfword immediate  
			latency_EX= 3-1; 	 
			imm_extended={ {6{imm10[9]}},imm10};
			RT[0+:16] = (~RA[0+:16]+1)+imm_extended;
			RT[16+:16]=(~RA[16+:16]+1)+imm_extended;
			RT[32+:16]=(~RA[32+:16]+1)+imm_extended;
			RT[48+:16]=(~RA[48+:16]+1)+imm_extended;
			RT[64+:16]=(~RA[64+:16]+1)+imm_extended;
			RT[80+:16]=(~RA[80+:16]+1)+imm_extended;
			RT[96+:16]=(~RA[96+:16]+1)+imm_extended;
			RT[112+:16]=(~RA[112+:16]+1)+imm_extended; 
		
	end 
	7'd11: //subtract from word
	begin 
		    latency_EX= 3-1; //subtract from word
			RT[0+:32] = (~RA[0+:32]+1)+RB[0+:32]; //bytes 0 and 3
			RT[32+:32]=(~RA[32+:32]+1)+RB[32+:32]; //bytes 4 and 7
			RT[64+:32]=(~RA[64+:32]+1)+RB[64+:32]; //bytes 8 and 11
			RT[96+:32]=(~RA[96+:32]+1)+RB[96+:32]; //bytes 12 and 15
			
		
		
	end   
	7'd12:
	begin 
			latency_EX= 3-1; //subtract from word immediate 
			imm_extended_32={ {22{imm10[9]}},imm10[9:0]};
			RT[0+:32] = (~RA[0+:32]+1)+imm_extended_32;
			RT[32+:32]=(~RA[32+:32]+1)+imm_extended_32;
			RT[64+:32]=(~RA[64+:32]+1)+imm_extended_32;
			RT[96+:32]=(~RA[96+:32]+1)+imm_extended_32; 
				
		
		
	end	  
	7'd13: begin //carry generate 
		RT=0;//set remaining bits to 0
		for(int j=0;j<16;j+=4) begin 
		temp_t[31:0]=(RA[j*8+:32]<<1)+(RB[j*8+:32]<<1);	
		RT[j*8+:32]=temp_t<<32;
		end  
		
		
		
	end 
	7'd14: begin //count leading zeros   
		latency_EX= 3-1; 
				for(int j=0;j<16;j+=4) begin 
					temp_32=32'd0;
					temp_u=RA[(j*8)+:32];
					for(int m=0;m<32;m+=1) begin 
						if(temp_u[m]==1) begin 
							break;  
							
						end	//end if
					else begin 
					temp_32=temp_32+1;	
						
					end //end else 
						
					end // end m loop
					
				RT[(j*8)+:32]=	temp_32;
				end// end for j loop
				
			end	 //end instr 
		7'd15: begin 	//and
			latency_EX= 3-1; 
		    RT[0+:32] = RA[0+:32]&RB[0+:32]; //bytes 0 and 3
			RT[32+:32]=RA[32+:32]&RB[32+:32]; //bytes 4 and 7
			RT[64+:32]=RA[64+:32]&RB[64+:32]; //bytes 8 and 11
			RT[96+:32]=RA[96+:32]&RB[96+:32]; //bytes 12 and 15
				
			
			
		end	 
		7'd16: begin //and with compliment
			latency_EX= 3-1; 
		    RT[0+:32] = RA[0+:32]&(~RB[0+:32]); //bytes 0 and 3
			RT[32+:32]=RA[32+:32]&(~RB[32+:32]); //bytes 4 and 7
			RT[64+:32]=RA[64+:32]&(~RB[64+:32]); //bytes 8 and 11
			RT[96+:32]=RA[96+:32]&(~RB[96+:32]); //bytes 12 and 15
				
	    end 
	   	7'd17: begin  //and halfword immediate 
			latency_EX= 3-1; 	 
			imm_extended={ {6{imm10[9]}},imm10};
			RT[0+:16] = RA[0+:16]&imm_extended;
			RT[16+:16]=RA[16+:16]&imm_extended;
			RT[32+:16]=RA[32+:16]&imm_extended;
			RT[48+:16]=RA[48+:16]&imm_extended;
			RT[64+:16]=RA[64+:16]&imm_extended;
			RT[80+:16]=RA[80+:16]&imm_extended;
			RT[96+:16]=RA[96+:16]&imm_extended;
			RT[112+:16]=RA[112+:16]&imm_extended;    
			   
	    end
		7'd18: begin //and word immediate
		    latency_EX= 3-1;   
	 		imm_extended_32={ {22{imm10[9]}},imm10[9:0]};
			RT[0+:32] = RA[0+:32]&imm_extended_32;
			RT[32+:32]=RA[32+:32]&imm_extended_32;
			RT[64+:32]=RA[64+:32]&imm_extended_32;
			RT[96+:32]=RA[96+:32]&imm_extended_32; 	
			
		end	  
		7'd19: begin //or 
			latency_EX= 3-1; 
		    RT[0+:32] = RA[0+:32]|RB[0+:32]; //bytes 0 and 3
			RT[32+:32]=RA[32+:32]|RB[32+:32]; //bytes 4 and 7
			RT[64+:32]=RA[64+:32]|RB[64+:32]; //bytes 8 and 11
			RT[96+:32]=RA[96+:32]|RB[96+:32]; //bytes 12 and 15
			
		end 
		7'd20: begin 	//or with complement 
			latency_EX= 3-1; 
		    	RT[0+:32] =RA[0+:32]|(~RB[0+:32]); //bytes 0 and 3
			RT[32+:32]=RA[32+:32]|(~RB[32+:32]); //bytes 4 and 7
			RT[64+:32]=RA[64+:32]|(~RB[64+:32]); //bytes 8 and 11
			RT[96+:32]=RA[96+:32]|(~RB[96+:32]); //bytes 12 and 15
				
			
		end 			
		7'd21: begin   //or halfword immediate 
					latency_EX= 3-1; 	 
			imm_extended={ {6{imm10}},imm10};
			RT[0+:16] = RA[0+:16]|imm_extended;
			RT[16+:16]=RA[16+:16]|imm_extended;
			RT[32+:16]=RA[32+:16]|imm_extended;
			RT[48+:16]=RA[48+:16]|imm_extended;
			RT[64+:16]=RA[64+:16]|imm_extended;
			RT[80+:16]=RA[80+:16]|imm_extended;
			RT[96+:16]=RA[96+:16]|imm_extended;
			RT[112+:16]=RA[112+:16]|imm_extended;    
			
		end 
		7'd22: begin    //or word immediate 
		    latency_EX= 3-1;   
	 		imm_extended_32={ {22{imm10[9]}},imm10[9:0]};
			RT[0+:32] = RA[0+:32]|imm_extended_32;
			RT[32+:32]=RA[32+:32]|imm_extended_32;
			RT[64+:32]=RA[64+:32]|imm_extended_32;
			RT[96+:32]=RA[96+:32]|imm_extended_32; 	
			
			
		end 
		7'd23: begin //exclusive or 
			latency_EX= 3-1; 
		    RT[0+:32] = RA[0+:32]^RB[0+:32]; //bytes 0 and 3
			RT[32+:32]=RA[32+:32]^RB[32+:32]; //bytes 4 and 7
			RT[64+:32]=RA[64+:32]^RB[64+:32]; //bytes 8 and 11
			RT[96+:32]=RA[96+:32]^RB[96+:32]; //bytes 12 and 15
			
		end  
		7'd24: begin    //exclusive or halfword immediate 
			latency_EX= 3-1; 	 
			imm_extended={ {6{imm10[9]}},imm10};
			RT[0+:16] = RA[0+:16]^imm_extended;
			RT[16+:16]=RA[16+:16]^imm_extended;
			RT[32+:16]=RA[32+:16]^imm_extended;
			RT[48+:16]=RA[48+:16]^imm_extended;
			RT[64+:16]=RA[64+:16]^imm_extended;
			RT[80+:16]=RA[80+:16]^imm_extended;
			RT[96+:16]=RA[96+:16]^imm_extended;
			RT[112+:16]=RA[112+:16]^imm_extended;  	
			
		end 
		7'd25: begin //exclusive or word immediate 
			 latency_EX= 3-1;   
	 		imm_extended_32={ {22{imm10[9]}},imm10[9:0]};
			RT[0+:32] = RA[0+:32]^imm_extended_32;
			RT[32+:32]=RA[32+:32]^imm_extended_32;
			RT[64+:32]=RA[64+:32]^imm_extended_32;
			RT[96+:32]=RA[96+:32]^imm_extended_32; 	
			
			
		end 
		7'd26: begin 	 //nand 
		   	latency_EX= 3-1; 
		    RT[0+:32] = ~(RA[0+:32]&RB[0+:32]); //bytes 0 and 3
			RT[32+:32]=~(RA[32+:32]&RB[32+:32]); //bytes 4 and 7
			RT[64+:32]=~(RA[64+:32]&RB[64+:32]); //bytes 8 and 11
			RT[96+:32]=~(RA[96+:32]&RB[96+:32]); //bytes 12 and 15
				
			
			
		end
		7'd76: begin 	 //nor 
			latency_EX= 3-1; 
		    RT[0+:32] = ~(RA[0+:32]|RB[0+:32]); //bytes 0 and 3
			RT[32+:32]=~(RA[32+:32]|RB[32+:32]); //bytes 4 and 7
			RT[64+:32]=~(RA[64+:32]|RB[64+:32]); //bytes 8 and 11
			RT[96+:32]=~(RA[96+:32]|RB[96+:32]); //bytes 12 and 15
			
		end 
		7'd28: begin 	//compare equal halfward
		latency_EX= 3-1;
		for(int j=0; j<16;j+=2) begin 
			if(RA[(j*8)+:16]==RB[(j*8)+:16]) begin 
				RT[(j*8)+:16]=11'hFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:16]=11'h00000;
			
		end 
			
		end 
			
			
		end	   
	7'd29: begin   //compare equal halfword immediate
		imm_extended={ {6{imm10[9]}},imm10};
	for(int j=0; j<16;j+=2) begin 
			if(RA[(j*8)+:16]==imm_extended) begin 
				RT[(j*8)+:16]=11'hFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:16]=11'h00000;
			
		end 
			
		end 
			
			
	end	
	7'd30: begin //compare equal word
			
	latency_EX= 3-1;
		for(int j=0; j<16;j+=4) begin 
			if(RA[(j*8)+:32]==RB[(j*8)+:32]) begin 
				RT[(j*8)+:32]=11'hFFFFFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:32]=11'h00000;
			
		end 
			
		end 
			
			
	end	  
	7'd31: begin  //compare equal word immediate
		latency_EX= 3-1;
		imm_extended_32={ {22{imm10[9]}},imm10};
	for(int j=0; j<16;j+=2) begin 
			if(RA[(j*8)+:32]==imm_extended_32) begin 
				RT[(j*8)+:32]=11'hFFFFFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:32]=11'h00000;
			
		end 
			
		end 
			
			
	end		
		
	 
	7'd32: begin 	  //compare greater than halfword
	latency_EX= 3-1;
		for(int j=0; j<16;j+=2) begin 
			if(RA[(j*8)+:16]>RB[(j*8)+:16]) begin 
				RT[(j*8)+:16]=11'hFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:16]=11'h00000;
			
		end 
			
		end 
			
			
		end	
		
	7'd33: begin //compare greater than halfword immediate
		latency_EX= 3-1;
		imm_extended={ {6{imm10[9]}},imm10};
	for(int j=0; j<16;j+=2) begin 
			if(RA[(j*8)+:16]>imm_extended) begin 
				RT[(j*8)+:16]=11'hFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:16]=11'h00000;
			
		end 
			
	end  
	
	end 
	 7'd34: begin //compare greater than word 
		latency_EX= 3-1;
		for(int j=0; j<16;j+=4) begin 
			if(RA[(j*8)+:32]>RB[(j*8)+:32]) begin 
				RT[(j*8)+:32]=11'hFFFFFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:32]=11'h00000;
			
		end 
			
		end 
			
			
	end	 
	7'd35: begin //compare greater than word immediate
		latency_EX= 3-1;
		imm_extended_32={ {22{imm10[9]}},imm10[9:0]};
	for(int j=0; j<16;j+=2) begin 
			if(RA[(j*8)+:32]>imm_extended_32) begin 
				RT[(j*8)+:32]=11'hFFFFFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:32]=11'h00000;
			
		end 
			
		end 
			
			
	end		
	7'd36: begin //compare logical greater than halfword

		latency_EX= 3-1;
		for(int j=0; j<16;j+=2) begin 
			if(unsigned_RA[(j*8)+:16]>unsigned_RB[(j*8)+:16]) begin 
				RT[(j*8)+:16]=11'hFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:16]=11'h00000;
			
		end 
			
		end 
			
			
		end	 
	7'd37: begin  //compare logical greater than halfword immediate 
	latency_EX= 3-1;
	imm_extended={ {6{imm10[9]}},imm10[9:0]}; 
	unsigned_imm_extended=unsigned'(imm_extended);
	for(int j=0; j<16;j+=2) begin 
			if(unsigned_RA[(j*8)+:16]>unsigned_imm_extended) begin 
				RT[(j*8)+:16]=11'hFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:16]=11'h00000;
			
		end 
			
	end  
	
	end 
	
	7'd38:  begin //compare logical greater than word
		latency_EX= 3-1;
		for(int j=0; j<16;j+=4) begin 
			if(unsigned_RA[(j*8)+:32]>unsigned_RB[(j*8)+:32]) begin 
				RT[(j*8)+:32]=11'hFFFFFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:32]=11'h00000;
			
		end 
			
		end 
			
			
	end	 
	7'd39: begin   //compare logical greater than word immediate 
			latency_EX= 3-1;
		imm_extended={ {6{imm10[9]}},imm10[9:0]};
		unsigned_imm_extended=unsigned'(imm_extended);
	for(int j=0; j<16;j+=2) begin 
			if(unsigned_RA[(j*8)+:16]>unsigned_imm_extended) begin 
				RT[(j*8)+:16]=11'hFFFF;
				
				
			end 
		else begin 
			RT[(j*8)+:16]=11'h00000;
			
		end 
			
	end  
	
	end  
	
	7'd40:begin //immediate load halfword
	latency_EX= 3-1;
	
	RT=imm16; 
		
	end 
	7'd41: begin //immediate load halfword upper
		latency_EX= 3-1;
			
		temp_t=imm16; //left shift by 16 to put in upper half
		RT=temp_t<<16; 
		
	end   
	7'd42: begin //imm load word
	latency_EX= 3-1;
	imm_extended_32={ {16{imm16[15]}},imm16};	
	RT=imm_extended_32; 
		
	end 
	7'd43: begin //immediate load address 
	latency_EX= 3-1;
	RT=imm18;
	RT[31:18]=0; //set rest of the bits to 0
		
	end 
	
	7'd44: begin //immediate or halfword lower
	latency_EX=3-1; 
	temp_t=imm16;
	temp_t[31:16]=0;  
	RT=RT|temp_t;
	
	
		
	end
	7'd45: begin //and byte immediate 
	temp_b=imm10 & 16'hFF;
	temp_bbbb[7:0]=temp_b;
	temp_bbbb[15:8]=temp_b;
	temp_bbbb[23:16]=temp_b;
	temp_bbbb[31:24]=temp_b;
	RT[0+:32]=RA[0+:24] &temp_bbbb;	  
	RT[32+:32]=RA[0+:24] &temp_bbbb;
	RT[64+:32]=RA[0+:24] &temp_bbbb;	 
	RT[96+:32]=RA[0+:24] &temp_bbbb;
		
	end 
	7'd46: begin 	//shift left halfword	
	for(int j=0;j<16;j+=2) begin 
   temp_s=RB[(j*8)+:16]&16'h1F; //halfword access +:16  
   temp_t=RA[(j*8)+:16];//halfword access +:16 
	for(int b=0;b<16;b++) begin 
   if((b+temp_s)<16) begin 
   temp_r[b]=temp_t[b+temp_s];

   end 
   else begin 
  temp_r[b]=0;

   end 


   end 

  RT[(j*8)+:16]=temp_r; //set 16 bits of register RT to r_temp  
  end 

   end 
		
   7'd47: begin //shift left halfword immediate 
	for(int j=0;j<16;j+=2) begin 
   imm_extended={ {11{imm7[6]}},imm7[6:0]};
   temp_s=imm_extended&16'h1F; //halfword access +:16  
   temp_t=RA[(j*8)+:16];//halfword access +:16 
	for(int b=0;b<16;b++) begin 
   if((b+temp_s)<16) begin 
   temp_r[b]=temp_t[b+temp_s];

   end 
   else begin 
  temp_r[b]=0;

   end 


   end    
     RT[(j*8)+:16]=temp_r; //set 16 bits of register RT to r_temp  
  end 

   end    
  7'd48: begin //shift left word
		for(int j=0;j<16;j+=4) begin 
   temp_s=RB[(j*8)+:32]&16'h3F; //halfword access +:16  
   temp_t=RA[(j*8)+:32];//halfword access +:16 
	for(int b=0;b<32;b++) begin 
   if((b+temp_s)<32) begin 
   temp_r[b]=temp_t[b+temp_s];

   end 
   else begin 
  temp_r[b]=0;

   end 


   end 

  RT[(j*8)+:32]=temp_r; //set 16 bits of register RT to r_temp  
  end 

   end   
	  
  7'd49: begin //shift left word immediate 
  	for(int j=0;j<32;j+=4) begin 
   imm_extended_32={ {25{imm7[6]}},imm7[6:0]};
   temp_s=imm_extended_32&16'h3F; //halfword access +:16  
   temp_t=RA[(j*8)+:32];//halfword access +:16 
	for(int b=0;b<32;b++) begin 
   if((b+temp_s)<32) begin 
   temp_r[b]=temp_t[b+temp_s];

   end 
   else begin 
  temp_r[b]=0;

   end 


   end    
     RT[(j*8)+:32]=temp_r; //set 16 bits of register RT to r_temp  
  end 

   end    
	  
  7'd86: begin 	  //Branch If Not Zero Word
	if(RT[0+:32]!=0) begin 
		 branch_flag=1; 
		 branch_PC=branch_PC_p2&32'hFFFFFFFC;
		
	end 
  else begin 
	branch_flag=0;   
	  
  end 
	  
	  
   end 
  7'd87: begin 	//branch if not zero halfword 
	if(RT[8+:16]!=0) begin 
		 branch_flag=1; 
		 branch_PC=branch_PC_p2&32'hFFFFFFFC;
		
	end 
  else begin 
	branch_flag=0;   
	  
  end 
	  
	  
   end 
	   
7'd90: begin  //branch if zero word 
	if(RT[0+:32]==0) begin 
		 branch_flag=1; 
		 branch_PC=branch_PC_p2&32'hFFFFFFFC;
		
	end 
  else begin 
	branch_flag=0;   
	  
  end 
	  
	  
   end 
/*7'd89: begin //branch if not zero halfword 
	if(RT[8+:16]!=0) begin 
		branch_flag=1;   
		branch_PC=branch_PC_p2&32'hFFFFFFFC;
		
		
	end 
  else begin 
	branch_flag=0;   
	  
  end 
	  
	  
   end */
  7'd91: begin 	//branch absolute
  branch_flag=1; 
	  
	  
end
7'd93: begin //branch relative
branch_flag=1;
branch_PC=branch_PC_p2; //removes mask from address
	
	
end 
7'd50: begin 	//rotate halfword 
	for(int j=0;j<16;j+=2) begin 
   temp_s=RB[(j*8)+:16]&16'hF; //halfword access +:16  
   temp_t=RA[(j*8)+:16];//halfword access +:16 
	for(int b=0;b<16;b++) begin 
   if((b+temp_s)<16) begin 
   temp_r[b]=temp_t[b+temp_s];

   end 
   else begin 
  temp_r[b]=temp_t[b+temp_s-16];

   end 


   end 

  RT[(j*8)+:16]=temp_r; //set 16 bits of register RT to r_temp  
  end 

   end  
7'd51: begin //rotate halfword immediate  
	for(int j=0;j<16;j+=2) begin 
   imm_extended={ {11{imm7[6]}},imm7[6:0]};
   temp_s=imm_extended&16'hF; //halfword access +:16  
   temp_t=RA[(j*8)+:16];//halfword access +:16 
	for(int b=0;b<16;b++) begin 
   if((b+temp_s)<16) begin 
   temp_r[b]=temp_t[b+temp_s];

   end 
   else begin 
  temp_r[b]=temp_t[b+temp_s-16];

   end 


   end    
     RT[(j*8)+:16]=temp_r; //set 16 bits of register RT to r_temp  
  end 

end  
7'd52: begin 	 //rotate word 
		for(int j=0;j<16;j+=4) begin 
   temp_s=RB[(j*8)+:32]&16'h1F; //word access +:16  
   temp_t=RA[(j*8)+:32];//word access +:16 
	for(int b=0;b<32;b++) begin 
   if((b+temp_s)<32) begin 
   temp_r[b]=temp_t[b+temp_s];

   end 
   else begin 
  temp_r[b]=temp_t[b+temp_s-32];

   end 


   end 

  RT[(j*8)+:32]=temp_r; //set 16 bits of register RT to r_temp  
  end 

end 
7'd53: begin //rotate word immediate 
	for(int j=0;j<32;j+=4) begin 
   imm_extended_32={ {25{imm7[6]}},imm7[6:0]};
   temp_s=imm_extended_32&16'h1F; //word access +:32  
   temp_t=RA[(j*8)+:32];//word access +:32 
	for(int b=0;b<32;b++) begin 
   if((b+temp_s)<32) begin 
   temp_r[b]=temp_t[b+temp_s];

   end 
   else begin 
  temp_r[b]=temp_t[b+temp_s-32];

   end 


   end    
     RT[(j*8)+:32]=temp_r; //set 16 bits of register RT to r_temp  
  end 

end 
7'd54: begin 			 //multiply op code 
		    RT[0+:32] = RA[0+:32]*RB[0+:32]; //bytes 0 and 3
			RT[32+:32]=RA[32+:32]*RB[32+:32]; //bytes 4 and 7
			RT[64+:32]=RA[64+:32]*RB[64+:32]; //bytes 8 and 11
			RT[96+:32]=RA[96+:32]*RB[96+:32]; //bytes 12 and 15
	
	
end   
7'd55: begin //multiply unsigned 
	        RT[0+:32] = unsigned_RA[0+:32]*unsigned_RB[0+:32]; //bytes 0 and 3
			RT[32+:32]=unsigned_RA[32+:32]*unsigned_RB[32+:32]; //bytes 4 and 7
			RT[64+:32]=unsigned_RA[64+:32]*unsigned_RB[64+:32]; //bytes 8 and 11
			RT[96+:32]=unsigned_RA[96+:32]*unsigned_RB[96+:32]; //bytes 12 and 15
	
end 
7'd56: begin  //multiply immediate 
            latency_EX= 3-1; //multiply word immediate	   
	 		imm_extended_32={ {22{imm10[9]}},imm10};
			RT[0+:32] = RA[0+:32]*imm_extended_32;
			RT[32+:32]=RA[32+:32]*imm_extended_32;
			RT[64+:32]=RA[64+:32]*imm_extended_32;
			RT[96+:32]=RA[96+:32]*imm_extended_32; 	
			
	
	
end 
7'd57: begin  //multiply unsigned immediate 
	        latency_EX= 3-1; //multiply word immediate	   
	 		imm_extended_32={ {22{imm10[9]}},imm10[9:0]};
			RT[0+:32] = unsigned_RA[0+:32]*unsigned'(imm_extended_32);
			RT[32+:32]=unsigned_RA[32+:32]*unsigned'(imm_extended_32);
			RT[64+:32]=unsigned_RA[64+:32]*unsigned'(imm_extended_32);
			RT[96+:32]=unsigned_RA[96+:32]*unsigned'(imm_extended_32); 	
	
	
end   
7'd58: begin //multiply and add
			temp_t = RA[0+:32]*RB[0+:32]; //bytes 0 and 3
			temp_t1=RA[32+:32]*RB[32+:32]; //bytes 4 and 7
			temp_t2=RA[64+:32]*RB[64+:32]; //bytes 8 and 11
			temp_t3=RA[96+:32]*RB[96+:32]; //bytes 12 and 15  
			RT[0+:32] = RC[0+:32]+temp_t;
			RT[32+:32]=RC[32+:32]+temp_t1;
			RT[64+:32]=RC[64+:32]+temp_t2;
			RT[96+:32]=RC[96+:32]+temp_t3; 	
	
	
	
	
end
7'd59: begin 	 //floating add 
RT=float_RA+float_RB;	
	
	
end  

7'd60: begin //floating subtract
RT=float_RA-float_RB;		
	
end  
7'd61:begin //floating multiply
RT=float_RA*float_RB;		
	
end 
7'd62:begin 		   //floating multiply and add 
RT=(float_RA*float_RB)+float_RC;	
	
end  

7'd63: begin //floating multiply and subtract 
RT=(float_RA*float_RB)-float_RC;	
	
	
end  
7'd64: begin //average bytes 
for(int j=0;j<16;j++) begin 
RT[(j*8)+:32]=(RA[(j*8)+:32]+RB[(j*8)+:32]+1)>>1;
	
	
end	
end 
7'd65: begin //counts ones in bytes 
for(int j=0;j<7;j++) begin 
	temp_c=0;
	temp_b=RA[(j*8)+:8];
	for(int m=0;m<7;m++) begin 
		if(temp_b==1) begin 
			
			temp_c=temp_c+1;
		end
	RT[(j*8)+:8]=temp_c;	
		
		
	end 
	
end 

end 
7'd66: begin //absolute differences of bytes 
	for(int j=0;j<16;j++) begin 
		if(unsigned_RB[(j*8)+:8]>unsigned_RA[(j*8)+:8]) begin 
			
		RT[(j*8)+:8]=unsigned_RB[(j*8)+:8]-unsigned_RA[(j*8)+:8];	
		end 
	else begin 
		RT[(j*8)+:8]=unsigned_RA[(j*8)+:8]-unsigned_RB[(j*8)+:8];	
		
	end 
		
	end 
	 

	
end	
7'd67: begin //sum bytes ito halfwords 
	RT[0+:16]=RB[0+:8]+RB[8+:8]+RB[16+:8]+RB[24+:8];  //bytes 0 and 1
	RT[16+:16]=RA[0+:8]+RA[8+:8]+RA[16+:8]+RA[24+:8];  //byes 2 and 3
	RT[32+:16]=RA[32+:8]+RA[40+:8]+RA[48+:8]+RA[56+:8];   //bytes 4 and 5
	RT[48+:16]=RB[32+:8]+RA[40+:8]+RA[48+:8]+RA[56+:8];	//bytes	 6 and 7
	RT[64+:16]=RB[64+:8]+RB[72+:8]+RB[80+:8]+RB[88+:8];//bytes 8 and 9 	  
	RT[80+:16]=RA[64+:8]+RA[72+:8]+RA[80+:8]+RA[88+:8];//bytes 10 and 11 
	RT[96+:16]=RB[96+:8]+RB[104+:8]+RB[112+:8]+RB[120+:8]; //bytes 12 and 13 
	RT[96+:16]=RA[96+:8]+RA[104+:8]+RA[112+:8]+RA[120+:8]; 	  //bytes 14 and 15
	
	
end   
7'd68: begin //compare equal byte
	for(int i=0;i<15;i++) begin 
		if(RA[(i*8)+:8]==RB[(i*8)+:8]) begin 
			RT[(i*8)+:8]=8'hFF;
			
		end 
	else begin 
		RT[(i*8)+:8]=0;
		
	end 
		
	end 
	
end
7'd69: begin //compare equal byte immediate 
for(int i=0;i<15;i++) begin 
		if(RA[(i*8)+:8]==imm10[2+:8]) begin 
			RT[(i*8)+:8]=8'hFF;
			
		end 
	else begin 
		RT[(i*8)+:8]=0;
		
	end 
		
end	
end 
7'd70: begin 	 //shift left quadword by bits 
	temp_s=RB[29+:3];
	for(int b=0;b<128;b++) begin 
		if((b+temp_s)<128) begin 
			temp_r[b]=RA[b+temp_s];
			
		end 
	else begin 
		temp_r[b]=0;
		
	end 
		
	end 
RT=temp_r;	
		
end 
7'd71: begin 		  //Shift Left Quadword by Bits Immediate
temp_s=imm7&7'h7;
for(int b=0;b<128;b++) begin 
		if((b+temp_s)<128) begin 
			temp_r[b]=RA[b+temp_s];
			
		end 
	else begin 
		temp_r[b]=0;
		
	end 
		
end
RT=temp_r;	
	
end 
7'd72: begin //shift left quadword by bytes 
	temp_s=RB[27+:5]; //bits 27-31 27,28,29,30,31 
for(int b=0;b<16;b++) begin 
	if(b+temp_s<16) begin 
		temp_r[(b*8)+:8]=RA[((b+temp_s)*8)+:8];
		
	end 
else begin 
	temp_r[(b*8)+:8]=0; 
end 
	
end 
RT=temp_r;	
	
end
7'd73: begin //shift left quadword by bytes immediate  	
	temp_s=imm7&7'h1F;
for(int b=0;b<16;b++) begin 
	if(b+temp_s<16) begin 
		temp_r[(b*8)+:8]=RA[((b+temp_s)*8)+:8];
		
	end 
else begin 
	temp_r[(b*8)+:8]=0; 
end 
	
end 
RT=temp_r;	
	
end	
7'd74: begin //shift left quadword by bits bit shift count 
	temp_s=RB[28:24]; //bits 24-28 24,25,26,27,28 
	for(int b=0; b<16;b++) begin 
		if((b+temp_s)<16) begin 
			temp_r[(b*8)+:8]=RA[((b+temp_s)*8)+:8];
			
		end   
	else begin 
		temp_r[(b*8)+:8]=0;
		
	end 
		
	end
	RT=temp_r;
end  
7'd75: begin 	  //rotate quadword by bytes 
temp_s=RB[31:28]; //28-31 28,29,30,31	
for(int b=0;b<16;b++) begin 
	if((b+temp_s)<16) begin 
		temp_r[(b*8)+:8]=RA[((b+temp_s)*8)+:8]; 
		
	end   
else begin 
temp_r[(b*8)+:8]=RA[((b+temp_s-16)*8)+:8]; 	
	
end 
	
end
RT=temp_r;
end 
7'd76: begin 	//rotate quadword by bytes immediate 
	 temp_s=imm7[14+:3]; //14,15,17
for(int b=0;b<16;b++) begin 
	if((b+temp_s)<16) begin 
		temp_r[(b*8)+:8]=RA[((b+temp_s)*8)+:8]; 
		
	end   
else begin 
temp_r[(b*8)+:8]=RA[((b+temp_s-16)*8)+:8]; 	
	
end 

end
RT=temp_r;
end 
7'd77: begin //rotate quadword by bits 
	for(int b=0;b<128;b++) begin 
		if((b+temp_s)<128) begin 
			temp_r[(b*8)+:8]=RA[((b+temp_s)*8)+:8];
		end  
		else begin 
temp_r[(b*8)+:8]=RA[((b+temp_s-128)*8)+:8]; 	
	
end 
	end  
RT=temp_r;	
end 
7'd78: begin //rotate quadword by bits immediate 
	temp_s=imm7[6:4]; 
	for(int b=0;b<128;b++) begin 
		if((b+temp_s)<128) begin 
			temp_r[(b*8)+:8]=RA[((b+temp_s)*8)+:8]; 
		end  
		else begin 
temp_r[(b*8)+:8]=RA[((b+temp_s-128)*8)+:8]; 	
	
end 
	end  
RT=temp_r;	
end 
7'd79: begin //gather bits from bytes 
	temp_k=0; 
	temp_s=0;
for(int j=7;j<128;j+=8) begin 
temp_s[temp_k]=RA[j];
temp_k=temp_k+1; 
	
end 
RT[0+:16]=0;
RT[16+:16]=temp_s; 
RT[(4*8)+:32]=0;
RT[(8*8)+:32]=0;
RT[(12*8)+:32]=0;
	
end 
7'd80: begin //gather bits from halfwords
	temp_k=0; 
	temp_s=0;
for(int j=15;j<128;j+=16) begin 
temp_s[temp_k]=RA[j];
temp_k=temp_k+1; 
	
end 
RT[0+:24]=0;
RT[24+:8]=temp_s; 
RT[(4*8)+:32]=0;
RT[(8*8)+:32]=0;
RT[(12*8)+:32]=0;
	
end 
7'd81: begin //gather bits from words 
	temp_k=0; 
	temp_s=0;
for(int j=31;j<128;j+=32) begin 
temp_s[temp_k]=RA[j];
temp_k=temp_k+1; 
	
end 
RT[0+:28]=0;
RT[28+:4]=temp_s; 
RT[(4*8)+:32]=0;
RT[(8*8)+:32]=0;
RT[(12*8)+:32]=0;
	
end
7'd82: begin  //load quadword d form
	//bits 0 to 3 of imm extended 32 is 0 
	//bits 4 to 13 should be 10 bits 
	//4,5,6,7,8,9,10,11,12,13 
	//18+14=32
	imm_extended_32[4:0]=0;
	imm_extended_32[13:4]=imm10;  
	
	imm_extended_32={{18{imm_extended_32[31]}},imm_extended_32};
	local_store_address=imm_extended_32+RA[0+:32]&32'hFFFFFFF0;
	RT=local_store_address;
	
end  
7'd83: begin //load quadword x form  

	local_store_address=(RB[0+:32]+RA[0+:32])&32'hFFFFFFF0;
	RT=local_store_address;
	
end 
7'd84: begin//store quadword d form  
    imm_extended_32={ imm10[9:0],{4{1'b0}}};
	imm_extended_32={{18{imm_extended_32[31]}},imm_extended_32};
	local_store_address=imm_extended_32+RA[0+:32]&32'hFFFFFFF0;
		
	
	
end 
7'd85: begin //store quadword x form 
	local_store_address=(RB[0+:32]+RA[0+:32])&32'hFFFFFFF0;
	
	
	
end 
endcase

end 								   
// ALU aluexecute(ALU_A,ALU_B,ALU_C,ALUControl,ALUResult,zero); // ALU Module
endmodule 



/*
module Execute_Testbench();
logic [127:0] readDataRA_EX; 
logic [127:0] readDataRB_EX;
logic [127:0] readDataRC_EX;
//where's register RT??????
logic [3:0] opcode_EX;
logic [127:0] result;
logic [10:0] opcode; 
logic [127:0] result_EX; //perhaps not needed, if we have  
assign opcode = 11'b00011001000; 
assign readDataRA_EX= 128'd543534534452345043;
assign readDataRB_EX= 128'd234234234545610253; 
Execute ex(readDataRA_EX,readDataRB_EX,readDataRC_EX,result,opcode,opcode_EX,result_EX);
endmodule
*/
