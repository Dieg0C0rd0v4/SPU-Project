
module shift3 (in, out);

input [10:0] in;
output [10:0] out;

assign out = in<<3; 


endmodule 
